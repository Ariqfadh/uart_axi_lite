
`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Reference Book: FPGA Prototyping By Verilog Examples Xilinx Spartan-3 Version
// Authored by: Dr. Pong P. Chu
// Published by: Wiley
//
// Adapted for the Basys 3 Artix-7 FPGA by David J. Marion
//
// Top Module for the Complete UART System
//
// Setup for 9600 Baud Rate
//
// For 9600 baud with 100MHz FPGA clock: 
// 9600 * 16 = 153,600
// 100 * 10^6 / 153,600 = ~651      (counter limit M)
// log2(651) = 10                   (counter bits N) 
//
// For 19,200 baud rate with a 100MHz FPGA clock signal:
// 19,200 * 16 = 307,200
// 100 * 10^6 / 307,200 = ~326      (counter limit M)
// log2(326) = 9                    (counter bits N)
//
// For 115,200 baud with 100MHz FPGA clock:
// 115,200 * 16 = 1,843,200
// 100 * 10^6 / 1,843,200 = ~52     (counter limit M)
// log2(52) = 6                     (counter bits N) 
//
// For 1500 baud with 100MHz FPGA clock:
// 1500 * 16 = 24,000
// 100 * 10^6 / 24,000 = ~4,167     (counter limit M)
// log2(4167) = 13                  (counter bits N) 
//
// Comments:
// - Many of the variable names have been changed for clarity
//////////////////////////////////////////////////////////////////////////////////

module uart_top
    #(
        parameter   DBITS = 8,
                    SB_TICK = 16,
                    FIFO_EXP = 2
    )
    (
        input  wire        clk_100MHz,
        input  wire        reset,
        input  wire        read_uart,
        input  wire        write_uart,
        input  wire        rx,
        input  wire [15:0] br_limit_in,  // Input baru untuk Baud Rate
        input  wire [DBITS-1:0] write_data,
        output wire        rx_full,
        output wire        rx_empty,
        output wire        tx,
        output wire [DBITS-1:0] read_data
    );
    
    wire tick;
    wire rx_done_tick;
    wire tx_done_tick;
    wire tx_empty;
    wire tx_fifo_not_empty;
    wire [DBITS-1:0] tx_fifo_out;
    wire [DBITS-1:0] rx_data_out;
    
    // Generator sekarang menerima input dinamis
    baud_rate_generator BAUD_RATE_GEN (
        .clk_100MHz(clk_100MHz), 
        .reset(reset),
        .M(br_limit_in), 
        .tick(tick)
    );
    
    uart_rx #(.DBITS(DBITS), .SB_TICK(SB_TICK)) UART_RX_UNIT (
        .clk_100MHz(clk_100MHz),
        .reset(reset),
        .rx(rx),
        .sample_tick(tick),
        .data_ready(rx_done_tick),
        .data_out(rx_data_out)
    );
    
    uart_tx #(.DBITS(DBITS), .SB_TICK(SB_TICK)) UART_TX_UNIT (
        .clk_100MHz(clk_100MHz),
        .reset(reset),
        .tx_start(tx_fifo_not_empty),
        .sample_tick(tick),
        .data_in(tx_fifo_out),
        .tx_done(tx_done_tick),
        .tx(tx)
    );
    
    fifo #(.DATA_SIZE(DBITS), .ADDR_SPACE_EXP(FIFO_EXP)) FIFO_RX_UNIT (
        .clk(clk_100MHz), .reset(reset),
        .write_to_fifo(rx_done_tick), .read_from_fifo(read_uart),
        .write_data_in(rx_data_out), .read_data_out(read_data),
        .empty(rx_empty), .full(rx_full)            
    );
       
    fifo #(.DATA_SIZE(DBITS), .ADDR_SPACE_EXP(FIFO_EXP)) FIFO_TX_UNIT (
        .clk(clk_100MHz), .reset(reset),
        .write_to_fifo(write_uart), .read_from_fifo(tx_done_tick),
        .write_data_in(write_data), .read_data_out(tx_fifo_out),
        .empty(tx_empty), .full()
    );
    
    assign tx_fifo_not_empty = ~tx_empty;
  
endmodule